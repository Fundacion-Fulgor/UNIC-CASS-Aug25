** sch_path: /foss/designs/UNIC-CASS-Aug25/sch/DLL/DLL_tb.sch
**.subckt DLL_tb
Vdd1 VDD GND 1.2
x1 VDD net1 va vc GND delay_variable
C4 vin2 GND 100f m=1
VIN3 net1 GND PULSE(0 1.2 0 5p 5p 1n 2n)
x9 VDD GND va vin2 large_delay_vto1p1
Vss1 VSS GND 0
x2 vin2 net2 net1 vdn phase_detector
x3 vup net3 vdn push_pull
**** begin user architecture code


.save v(vin1) v(vin2)  v(vc) v(vdn) v(vup)



.tran 10p 10n
.save all
*.ic v(vout) = 0
.control
run
plot v(vin1) v(vin2)
plot v(vc)
plot v(vup) v(vdn)


*plot v(vin2)

*plot v(vout)
*meas tran teval WHEN v(vout) = 0.63
*let res_val = 1000
*let cap_val = teval/res_val
*print cap_val
.endc



.lib cornerMOSlv.lib mos_tt
.include /foss/pdks/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice

**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/UNIC-CASS-Aug25/sym/delay_variable/delay_variable.sym # of pins=5
** sym_path: /foss/designs/UNIC-CASS-Aug25/sym/delay_variable/delay_variable.sym
** sch_path: /foss/designs/UNIC-CASS-Aug25/sym/delay_variable/delay_variable.sch
.subckt delay_variable VDD_D VIN_D VOUT_D VCONT_D VSS_D
*.iopin VSS_D
*.iopin VDD_D
*.opin VOUT_D
*.ipin VCONT_D
*.ipin VIN_D
XM3 net4 VCONT_D net2 net2 sg13_lv_nmos w=1u l=0.13u ng=1 m=1
XM5 net3 VCONT_D net2 net2 sg13_lv_nmos w=2u l=2u ng=1 m=1
XM4 net4 net4 VDD_D VDD_D sg13_lv_pmos w=2.24*1u l=0.13u ng=1 m=1
XM6 net1 net4 VDD_D VDD_D sg13_lv_pmos w=4*1u l=2u ng=1 m=1
XM7 VOUT_D VIN_D net1 VDD_D sg13_lv_pmos w=4*5u l=2u ng=4 m=1
XM8 VOUT_D VIN_D net3 net2 sg13_lv_nmos w=5u l=3u ng=1 m=1
.ends


* expanding   symbol:  /foss/designs/UNIC-CASS-Aug25/sym/large_delay_vto1p1/large_delay_vto1p1.sym # of pins=4
** sym_path: /foss/designs/UNIC-CASS-Aug25/sym/large_delay_vto1p1/large_delay_vto1p1.sym
** sch_path: /foss/designs/UNIC-CASS-Aug25/sym/large_delay_vto1p1/large_delay_vto1p1.sch
.subckt large_delay_vto1p1 VCC VSS VIN VOUT
*.iopin VIN
*.iopin VOUT
*.iopin VCC
*.iopin VSS
x1 VIN VCC VSS VOUT sg13g2_dlygate4sd1_1
x2 VIN VCC VSS VOUT sg13g2_dlygate4sd1_1
x3 VIN VCC VSS VOUT sg13g2_dlygate4sd1_1
x4 VIN VCC VSS VOUT sg13g2_dlygate4sd1_1
.ends


* expanding   symbol:  /foss/designs/UNIC-CASS-Aug25/sym/phase_detector/phase_detector.sym # of pins=4
** sym_path: /foss/designs/UNIC-CASS-Aug25/sym/phase_detector/phase_detector.sym
** sch_path: /foss/designs/UNIC-CASS-Aug25/sym/phase_detector/phase_detector.sch
.subckt phase_detector CK_IN UP CK_REF DN
*.opin UP
*.opin DN
*.ipin CK_IN
*.ipin CK_REF
XM7 net2 CK_IN VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM8 net1 CK_IN VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM9 net2 CK_REF net1 net1 sg13_lv_nmos w=2u l=5u ng=5 m=1
XM10 net2 DN net1 VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM11 net1 CK_IN VSS VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM6 net7 net6 VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM12 net7 CK_IN net8 net9 sg13_lv_nmos w=2u l=5u ng=5 m=1
XM13 net8 net6 net9 net9 sg13_lv_nmos w=2u l=5u ng=5 m=1
XM14 net8 net6 VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM1 net11 CK_IN VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM2 net10 CK_IN VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM3 net11 CK_REF net10 net10 sg13_lv_nmos w=2u l=5u ng=5 m=1
XM4 net11 UP net10 VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM5 net10 CK_IN VSS VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM15 net14 net13 VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM16 net14 CK_REF net15 VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM17 net15 net13 VSS VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM18 net15 net13 VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
x1 VDD net2 net3 net5 inv_1_manual
x7 VDD net3 net6 net4 inv_1_manual
x2 VDD net11 net12 VSS inv_1_manual
x8 VDD net12 net13 VSS inv_1_manual
x3 VDD net14 DN VSS inv_1_manual
x4 VDD net7 UP net9 inv_1_manual
.ends


* expanding   symbol:  /foss/designs/UNIC-CASS-Aug25/sym/push_pull/push_pull.sym # of pins=3
** sym_path: /foss/designs/UNIC-CASS-Aug25/sym/push_pull/push_pull.sym
** sch_path: /foss/designs/UNIC-CASS-Aug25/sym/push_pull/push_pull.sch
.subckt push_pull UP_IN VC DN_IN
*.ipin DN_IN
*.ipin UP_IN
*.opin VC
XM1 net1 DN_IN net2 VSS sg13_lv_nmos w=0.3u l=0.45u ng=1 m=1
XM7 net1 net1 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM2 net7 DNB net2 VSS sg13_lv_nmos w=0.3u l=0.45u ng=1 m=1
XM3 net2 VDD VSS VSS sg13_lv_nmos w=0.3u l=0.45u ng=1 m=1
XM4 net1 net1 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM5 net5 net7 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM6 net4 UPB net3 VSS sg13_lv_nmos w=0.3u l=0.45u ng=1 m=1
XM8 net6 net4 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM9 VC UP_IN net3 VSS sg13_lv_nmos w=0.3u l=0.45u ng=1 m=1
XM10 net3 VDD VSS VSS sg13_lv_nmos w=0.3u l=0.45u ng=1 m=1
XM11 VC net1 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM12 VC net1 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM13 net6 net4 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM14 net5 net7 VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
x1 VDD DN_IN DNB VSS inv_1_manual
x2 VDD UP_IN UPB VSS inv_1_manual
C1 VC VSS 10f m=1
.ends


* expanding   symbol:  /foss/designs/UNIC-CASS-Aug25/sym/inv_1_manual/inv_1_manual.sym # of pins=4
** sym_path: /foss/designs/UNIC-CASS-Aug25/sym/inv_1_manual/inv_1_manual.sym
** sch_path: /foss/designs/UNIC-CASS-Aug25/sym/inv_1_manual/inv_1_manual.sch
.subckt inv_1_manual VDD_D A Y VSS_D
*.iopin VDD_D
*.iopin VSS_D
*.iopin A
*.iopin Y
XM1 Y A VSS_D VSS_D sg13_lv_nmos w=10u l=0.13u ng=1 m=1
XM2 Y A VDD_D VDD_D sg13_lv_pmos w=10u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
