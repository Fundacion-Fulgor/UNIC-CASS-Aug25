** sch_path: /home/designer/UNIC-CASS-Aug25/Custom_std_cells/and_custom.sch
**.subckt and_custom VDD A OUT B VSS
*.ipin A
*.iopin VDD
*.opin OUT
*.iopin VSS
*.ipin B
x2 VDD OUT net1 VSS inv
x1 VDD net2 A B VSS nand_custom
**.ends

* expanding   symbol:  inv.sym # of pins=4
** sym_path: /home/designer/UNIC-CASS-Aug25/Custom_std_cells/inv.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/Custom_std_cells/inv.sch
.subckt inv VDD VOUT VIN VSS
*.iopin VDD
*.iopin VSS
*.opin VOUT
*.ipin VIN
XM2 VOUT VIN VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=2
XM1 VOUT VIN VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  nand_custom.sym # of pins=5
** sym_path: /home/designer/UNIC-CASS-Aug25/Custom_std_cells/nand_custom.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/Custom_std_cells/nand_custom.sch
.subckt nand_custom VDD OUT A B VSS
*.iopin A
*.iopin B
*.iopin VDD
*.iopin VSS
*.iopin OUT
XM1 OUT A net1 VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 OUT A VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 net1 B VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 OUT B VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends

.end
