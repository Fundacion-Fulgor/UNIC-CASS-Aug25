** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/tb_Circuit_stdcells.sch
**.subckt tb_Circuit_stdcells
C1 net1 avss 1p m=1
C2 net4 avss 1p m=1
C3 net2 avss 1p m=1
C4 net3 avss 1p m=1
V1 avss GND DC{vss}
V2 avdd avss DC{vdd}
V3 vs3 avss DC{a} PULSE(0 {vdd} 0.0 1p 1p {2*Tclk} {4*Tclk}) AC 0
V4 vs4 avss DC={vdd*c+1.2*d} PULSE(0 {vdd} 0.0 1p 1p {Tclk} {2*Tclk}) AC 0
x1 vs4 vs3 vo_s1t vo_s2t vo_s3t avdd vo_s4t avss Circuit_stdcells
x2 avdd vo_s1t net1 avss inv_prtt
x3 avdd vo_s2t net4 avss inv_prtt
x4 avdd vo_s3t net2 avss inv_prtt
x5 avdd vo_s4t net3 avss inv_prtt
B1 net5 net6 I = 'pwl(V(plus,minus),0,0, 1,10m, 2, 100m)' m=1
**** begin user architecture code



* Circuit Parameters
.param vdd = 1.2
.param vss = 0.0
.csparam VDD={vdd}
.csparam VSS={vss}
.param a=0
.param b=0
.param c=0
.param d=0
.param Tclk = 500n
.param a=0
.param b=0
.options TEMP = 65.0

* Include Models
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ


*.lib cornerMOSlv.lib mos_tt
*.lib cornerMOShv.lib mos_tt
*.lib cornerHBT.lib hbt_typ
*.lib cornerRES.lib res_typ
*.lib cornerCAP.lib cap_typ

* OP Parameters & Singals to save
.save all

*Simulations
.control
	tran 0.02u 10u
	setplot tran1
	plot v(vs4)+(5*2) v(vs3)+(4*2) v(vo_s1t)+(3*2) v(vo_s2t)+(2*2) v(vo_s3t)+2 v(vo_s4t) ylimit 0 12
	reset
	*dc @V3[a] 0 1.2 0.01
	let start_a=0
	let stop_a=1.2
	let delta_a=0.01
	let a_act=start_a
	while a_act le stop_a
		alterparam a = a_act
		reset
		run
		let a_act=a_act+delta_a
	end
	setplot dc1
	plot vo_s3t vs4 vs3 ylabel vout xlabel vin xlimit 0.55 0.65
	reset
	alter
	dc V3 0 1.2 0.01
	setplot dc2
	plot v(vo_s3t) v(vo_s2t) v(vs3) v(vs4) xlimit 0.55 0.65
	reset
	dc V3 0 1.2 0.01
	setplot dc3
	plot v(vo_s3t) v(vo_s2t) v(vs3) v(vs4) xlimit 0.55 0.65
.endc
.end

**** end user architecture code
**.ends

* expanding   symbol:  /home/designer/UNIC-CASS-Aug25/BinarytoThermo/Circuit_stdcells.sym # of pins=8
** sym_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/Circuit_stdcells.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/Circuit_stdcells.sch
.subckt Circuit_stdcells s4 s3 s1t s2t s3t vdd s4t vss
*.iopin s4
*.iopin s3
*.iopin s1t
*.iopin s2t
*.iopin s3t
*.iopin s4t
*.iopin vdd
*.iopin vss
x3 vdd s3t net1 net2 vss nand_prtt
x1 vdd net1 s1t net2 vss nor_prtt
x2 vdd s4 net1 vss inv_prtt
x4 vdd net2 s2t vss inv_prtt
x5 vdd s3 net2 vss inv_prtt
x6 vdd vss s4t vss inv_prtt
.ends


* expanding   symbol:  /home/designer/UNIC-CASS-Aug25/BinarytoThermo/inv_prtt.sym # of pins=4
** sym_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/inv_prtt.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/inv_prtt.sch
.subckt inv_prtt vdd in out vss
*.iopin in
*.iopin out
*.iopin vdd
*.iopin vss
XM1 out in vss vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 out in vdd vdd sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nand_prtt.sym # of pins=5
** sym_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nand_prtt.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nand_prtt.sch
.subckt nand_prtt vdd out A B vss
*.iopin A
*.iopin B
*.iopin vdd
*.iopin vss
*.iopin out
XM1 out A net1 vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 out A vdd vdd sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 net1 B vss vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 out B vdd vdd sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nor_prtt.sym # of pins=5
** sym_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nor_prtt.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nor_prtt.sch
.subckt nor_prtt vdd A out B vss
*.iopin vdd
*.iopin vss
*.iopin A
*.iopin B
*.iopin out
XM1 out B vss vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 out B net1 vdd sg13_lv_pmos w=0.45u l=0.13u ng=1 m=1
XM3 out A vss vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 net1 A vdd vdd sg13_lv_pmos w=0.45u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
