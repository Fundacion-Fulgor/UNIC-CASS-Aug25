** sch_path: /home/designer/shared/UNIC-CASS-Aug25/tb_delaycell.sch
**.subckt tb_delaycell
Vin1 in GND dc 0 ac 0 pulse(0, 1.2, 0, 25p, 25p, 250p, 500p )
Vdd1 net1 GND 1.2
C2 net3 net4 1f m=1
VCONT net2 net5 dc {VCONT}
x1 net1 in out net2 GND variable_delay
**** begin user architecture code

.lib cornerMOSlv.lib mos_tt



.param temp=27
.Param VCONT=0.9
.control
  save all
  step param VCONT 0.40 0.90 0.05   ; barrido 0.40→0.90 V en pasos de 50 mV
   *Vcont vcont 0 PWL(0n 0.40 10n 0.90)
  tran 1p 3n
  *meas tran tdelay TRIG v(in) VAL=0.9 FALL=1 TARG v(out) VAL=0.9 RISE=1
  write tran_logic_not.raw
.endc
.end


**** end user architecture code
**.ends

* expanding   symbol:  variable_delay.sym # of pins=5
** sym_path: /home/designer/shared/UNIC-CASS-Aug25/variable_delay.sym
** sch_path: /home/designer/shared/UNIC-CASS-Aug25/variable_delay.sch
.subckt variable_delay VDD VIN VOUT VCONT VSS
*.iopin VSS
*.iopin VDD
*.ipin VIN
*.opin VOUT
*.ipin VCONT
XM5 net2 VCONT VSS VSS sg13_lv_nmos w=5u l=0.13u ng=1 m=1
XM6 net1 net3 VDD VDD sg13_lv_pmos w=5u l=0.13u ng=1 m=1
XM2 VOUT VIN net1 VDD sg13_lv_pmos w=0.88u l=0.13u ng=4 m=1
XM1 VOUT VIN net2 VSS sg13_lv_nmos w=0.4u l=0.13u ng=1 m=1
x1 VDD VCONT net3 VSS inv_1_manual
.ends


* expanding   symbol:  /home/designer/shared/UNIC-CASS-Aug25/others/inv_1_manual.sym # of pins=4
** sym_path: /home/designer/shared/UNIC-CASS-Aug25/others/inv_1_manual.sym
** sch_path: /home/designer/shared/UNIC-CASS-Aug25/others/inv_1_manual.sch
.subckt inv_1_manual VDD_D A Y VSS_D
*.iopin VDD_D
*.iopin VSS_D
*.iopin A
*.iopin Y
XM1 Y A VSS_D VSS_D sg13_lv_nmos w=10u l=0.13u ng=1 m=1
XM2 Y A VDD_D VDD_D sg13_lv_pmos w=10u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
