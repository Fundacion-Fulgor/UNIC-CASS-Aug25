** sch_path: /home/designer/shared/UNIC-CASS-Aug25/phase_detector.sch
**.subckt phase_detector CK_IN UP CK_REF DN
*.opin UP
*.opin DN
*.ipin CK_IN
*.ipin CK_REF
XM7 net2 CK_IN VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM8 net1 CK_IN VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM9 net2 CK_REF net1 net1 sg13_lv_nmos w=2u l=5u ng=5 m=1
XM10 net2 DN net1 VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM11 net1 CK_IN VSS VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM6 net7 net6 VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM12 net7 CK_IN net8 net9 sg13_lv_nmos w=2u l=5u ng=5 m=1
XM13 net8 net6 net9 net9 sg13_lv_nmos w=2u l=5u ng=5 m=1
XM14 net8 net6 VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM1 net11 CK_IN VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM2 net10 CK_IN VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM3 net11 CK_REF net10 net10 sg13_lv_nmos w=2u l=5u ng=5 m=1
XM4 net11 UP net10 VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM5 net10 CK_IN VSS VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM15 net14 net13 VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
XM16 net14 CK_REF net15 VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM17 net15 net13 VSS VSS sg13_lv_nmos w=2u l=5u ng=5 m=1
XM18 net15 net13 VDD VDD sg13_lv_pmos w=5u l=4u ng=1 m=1
x1 VDD net11 net12 VSS inv_1_manual
x2 VDD net12 net13 VSS inv_1_manual
x3 VDD net14 DN VSS inv_1_manual
x4 VDD net7 UP net9 inv_1_manual
x5 VDD net3 net6 net4 inv_1_manual
x6 VDD net2 net3 net5 inv_1_manual
**.ends

* expanding   symbol:  /home/designer/shared/UNIC-CASS-Aug25/others/inv_1_manual.sym # of pins=4
** sym_path: /home/designer/shared/UNIC-CASS-Aug25/others/inv_1_manual.sym
** sch_path: /home/designer/shared/UNIC-CASS-Aug25/others/inv_1_manual.sch
.subckt inv_1_manual VDD_D A Y VSS_D
*.iopin VDD_D
*.iopin VSS_D
*.iopin A
*.iopin Y
XM1 Y A VSS_D VSS_D sg13_lv_nmos w=10u l=0.13u ng=1 m=1
XM2 Y A VDD_D VDD_D sg13_lv_pmos w=10u l=0.13u ng=1 m=1
.ends

.end
