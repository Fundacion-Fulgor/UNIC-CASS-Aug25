** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/tb_Circuit_stdcells_tran.sch
**.subckt tb_Circuit_stdcells_tran
C1 net1 avss 1p m=1
C2 net4 avss 1p m=1
C3 net2 avss 1p m=1
C4 net3 avss 1p m=1
V1 avss GND DC{vss}
V2 avdd avss DC{vdd}
V4 vs3 avss PULSE({a*1.2} {b*1.2} 250PS 2PS 2PS 500PS) DC 0
x1 vs4 vs3 vo_s1t vo_s2t vo_s3t avdd vo_s4t avss Circuit_stdcells
x2 avdd vo_s1t net1 avss inv_prtt
x3 avdd vo_s2t net4 avss inv_prtt
x4 avdd vo_s3t net2 avss inv_prtt
x5 avdd vo_s4t net3 avss inv_prtt
V7 vs4 avss PULSE({c*1.2} {d*1.2} 250PS 2PS 2PS 500PS)
**** begin user architecture code



* Circuit Parameters
.param vdd = 1.2
.param vss = 0.0
.param a=0
.param b=0
.param c=0
.param d=1
.param Tclk = 500P
.options TEMP = 65.0

* Include Models
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerMOShv.lib mos_tt
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerHBT.lib hbt_typ
.lib /opt/pdks/ihp-sg13g2/libs.tech/ngspice/models/cornerRES.lib res_typ


* OP Parameters & Singals to save
.save all

*Simulations
.control
set output_path = tb_termopi_tran/
	* Desde (s3,s4)=00 a 01
	tran 0.2PS 750PS
	setplot tran1
	plot vs3 vs4 vo_s3t ylabel vout xlabel vin
	set filetype = ascii
	write {$output_path}tran00to01.raw V(vo_s3t) V(vs3) V(vs4)
	* Desde (s3,s4)=00 a 10
	alterparam d=0
	alterparam b=1
	reset
	tran 0.2PS 750PS
	setplot tran2
	plot vs3 vs4 vo_s2t vo_s3t ylabel vout xlabel vin
	set filetype = ascii
	write {$output_path}tran00to10.raw V(vo_s2t) V(vo_s3t) V(vs3) V(vs4)
	* Desde (s3,s4)=00 a 11
	alterparam d = 1
	reset
	tran 0.2PS 750PS
	setplot tran3
	plot vs3 vs4 vo_s1t vo_s2t vo_s3t ylabel vout xlabel vin
	set filetype = ascii
	write {$output_path}tran00to11.raw V(vo_s1t) V(vo_s2t) V(vo_s3t) V(vs3) V(vs4)
	* Desde (s3,s4)=01 a 10
	alterparam c=1
	alterparam d=0
	reset
	tran 0.2PS 750PS
	setplot tran4
	plot vs3 vs4 vo_s2t ylabel vout xlabel vin
	set filetype = ascii
	write {$output_path}tran01to10.raw V(vo_s2t) V(vs3) V(vs4)
	* Desde (s3,s4)=01 a 11
	alterparam a=0
	alterparam b=1
	alterparam d=1
	reset
	tran 0.2PS 750PS
	setplot tran5
	plot vs3 vs4 vo_s1t vo_s2t ylabel vout xlabel vin
	set filetype = ascii
	write {$output_path}tran01to11.raw V(vo_s1t) V(vo_s2t) V(vs3) V(vs4)
	* Desde (s3,s4)=10 a 11
	alterparam a=1
	alterparam c=0
	alterparam d=1
	reset
	tran 0.2PS 750PS
	setplot tran6
	plot vs3 vs4 vo_s1t ylabel vout xlabel vin ylimit 0 1.2
	set filetype = ascii
	write {$output_path}tran10to11.raw V(vo_s1t) V(vs3) V(vs4)
.endc
.end

**** end user architecture code
**.ends

* expanding   symbol:  /home/designer/UNIC-CASS-Aug25/BinarytoThermo/Circuit_stdcells.sym # of pins=8
** sym_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/Circuit_stdcells.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/Circuit_stdcells.sch
.subckt Circuit_stdcells s4 s3 s1t s2t s3t vdd s4t vss
*.iopin s4
*.iopin s3
*.iopin s1t
*.iopin s2t
*.iopin s3t
*.iopin s4t
*.iopin vdd
*.iopin vss
x3 vdd s3t net1 net2 vss nand_prtt
x1 vdd net1 s1t net2 vss nor_prtt
x2 vdd s4 net1 vss inv_prtt
x4 vdd net2 s2t vss inv_prtt
x5 vdd s3 net2 vss inv_prtt
x6 vdd vss s4t vss inv_prtt
.ends


* expanding   symbol:  /home/designer/UNIC-CASS-Aug25/BinarytoThermo/inv_prtt.sym # of pins=4
** sym_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/inv_prtt.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/inv_prtt.sch
.subckt inv_prtt vdd in out vss
*.iopin in
*.iopin out
*.iopin vdd
*.iopin vss
XM1 out in vss vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 out in vdd vdd sg13_lv_pmos w=0.3u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nand_prtt.sym # of pins=5
** sym_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nand_prtt.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nand_prtt.sch
.subckt nand_prtt vdd out A B vss
*.iopin A
*.iopin B
*.iopin vdd
*.iopin vss
*.iopin out
XM1 out A net1 vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 out A vdd vdd sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
XM3 net1 B vss vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 out B vdd vdd sg13_lv_pmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nor_prtt.sym # of pins=5
** sym_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nor_prtt.sym
** sch_path: /home/designer/UNIC-CASS-Aug25/BinarytoThermo/nor_prtt.sch
.subckt nor_prtt vdd A out B vss
*.iopin vdd
*.iopin vss
*.iopin A
*.iopin B
*.iopin out
XM1 out B vss vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 out B net1 vdd sg13_lv_pmos w=0.45u l=0.13u ng=1 m=1
XM3 out A vss vss sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM4 net1 A vdd vdd sg13_lv_pmos w=0.45u l=0.13u ng=1 m=1
.ends

.GLOBAL GND
.end
