** sch_path: /home/designer/shared/martin.sch
.subckt martin

M9 VN2 VN2 VDD VDD sg13_lv_pmos w=0.52u l=0.26u ng=1 m=1
M6 net1 VN2 VDD VDD sg13_lv_pmos w=6u l=0.26u ng=1 m=1
M2 VOUT VIN net1 VDD sg13_lv_pmos w=8u l=0.26u ng=1 m=1
M8 VN2 Vctrl VSS VSS sg13_lv_nmos w=0.26u l=0.26u ng=1 m=1
M7 net2 Vctrl VSS VSS sg13_lv_nmos w=3.0u l=0.26u ng=1 m=1
M1 VOUT VIN net2 VSS sg13_lv_nmos w=4u l=0.26u ng=1 m=1
VDD VDD GND 1.2
VSS1 VSS GND 0
VIN1 VIN VSS PULSE(0 1.2 0 0.1p 0.1p 71.5p 143p)
VDD1 Vctrl GND 1.2
.ends
.GLOBAL GND
