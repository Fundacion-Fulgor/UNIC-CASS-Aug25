** sch_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/UNIC-CASS-Aug25/Differential_OTA_Telescopic_IHP/OTA_Telescopic_TB2_STB.sch
**.subckt OTA_Telescopic_TB2_STB
V7 vcm1 GND 1.25
V1 VDD GND 1.98
V2 VREF GND 0.9
C1 Vout2 GND 500f m=1
C2 Vout1 GND 500f m=1
R5 net1 vcm1 3k m=1
R6 net2 vcm1 3k m=1
I1 VDD net3 105u
x1 VDD vf1 Vout2 Vout1 vcm1 vcm1 GND net3 OTA_Telescopic_core_v2
x2 VDD VREF Vout1 Vout2 net4 vr1 GND OTA_Telescopic_CMFB2
I2 net4 GND 105u
R1 Vout2 net2 6.72k m=1
R2 Vout1 net1 6.72k m=1
Vtest1 vr1 vf1 dc 0 ac 1
V3 vcm2 GND 1.25
C3 V2 GND 500f m=1
C4 V1 GND 500f m=1
R7 net7 vcm2 3k m=1
R8 net8 vcm2 3k m=1
I3 VDD net5 105u
x3 VDD cmfb1 V2 V1 vcm2 vcm2 GND net5 OTA_Telescopic_core_v2
x4 VDD VREF V1 V2 net6 net24 GND OTA_Telescopic_CMFB2
I4 net6 GND 105u
R9 V2 net8 6.72k m=1
R10 V1 net7 6.72k m=1
Vif1 net9 cmfb1 0
.save i(vif1)
Vir1 net24 net9 0
.save i(vir1)
Itest1 GND net9 dc 0 ac 1
V4 net10 GND 1.2
C5 Vout22 GND 500f m=1
C6 Vout11 GND 500f m=1
I5 VDD net13 100u
x5 VDD vmeas1 Vout22 Vout11 net10 net10 GND net13 OTA_Telescopic_core_v2
x6 VDD VREF Vout22 Vout11 net14 net15 GND OTA_Telescopic_CMFB2
I6 net14 GND 100u
V5 net16 GND 1.2
C7 V22 GND 500f m=1
C8 V11 GND 500f m=1
I7 VDD net19 100u
x7 VDD vmeas2 V22 V11 net16 net16 GND net19 OTA_Telescopic_core_v2
x8 VDD VREF V22 V11 net20 net21 GND OTA_Telescopic_CMFB2
I8 net20 GND 100u
R21 net10 net11 10G m=1
R22 net10 net12 10G m=1
R23 net16 net17 10G m=1
R24 net16 net18 10G m=1
Vtest3 vmeas1 net22 dc 0 ac 1
Vimeas1 net15 net22 0
.save i(vimeas1)
Vtest2 vmeas2 net23 dc 0 ac 0
Vimeas2 net21 net23 0
.save i(vimeas2)
Itest2 GND vmeas1 dc 0 ac 0
Itest3 GND vmeas2 dc 0 ac 1
R3 vcm1 net1 10G m=1
R4 vcm1 net2 10G m=1
R11 vcm2 net7 10G m=1
R12 vcm2 net8 10G m=1
R13 net12 net10 3k m=1
R14 net11 net10 3k m=1
R15 net17 net16 3k m=1
R16 net18 net16 3k m=1
R17 Vout11 net11 6.72k m=1
R18 Vout22 net12 6.72k m=1
R19 V11 net17 6.72k m=1
R20 V22 net18 6.72k m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib cornerMOSlv.lib mos_ff
.temp 0



.op

.save all
*OTA
.save @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
.save @m.x1.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]

.save @m.x1.xm9.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x1.xm9.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x1.xm10.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x1.xm10.msky130_fd_pr__pfet_01v8_lvt[gm]

.save @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[id]

.save @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[vdssat]


.save @m.x1.xm13.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm14.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm15.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x1.xm16.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm17.msky130_fd_pr__nfet_01v8_lvt[id]

.save @m.x1.xm18.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x1.xm19.msky130_fd_pr__nfet_01v8_lvt[id]

*CMFB
.save @m.x2.xm0.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm1.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm1.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm2.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm2.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm3.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm4.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm4.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm5.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm6.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm6.msky130_fd_pr__pfet_01v8_lvt[gm]

.save @m.x2.xm7.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x2.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]
.save @m.x2.xm8.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x2.xm8.msky130_fd_pr__nfet_01v8_lvt[gm]



.control

let vdssat_M1 = @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[vdsat]
let vdssat_M3 = @m.x1.xm3.msky130_fd_pr__nfet_01v8_lvt[vdsat]
let vdssat_M5 = @m.x1.xm5.msky130_fd_pr__pfet_01v8_lvt[vdsat]
let vdssat_M7 = @m.x1.xm7.msky130_fd_pr__pfet_01v8_lvt[vdsat]
let vdssat_M0 = @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[vdsat]

let vdssat_M9 = @m.x1.xm9.msky130_fd_pr__pfet_01v8_lvt[vdsat]
let vdssat_M11 = @m.x1.xm11.msky130_fd_pr__nfet_01v8_lvt[vdsat]

print vdssat_M1
print vdssat_M3
print vdssat_M5
print vdssat_M7
print vdssat_M0
print vdssat_M9
print vdssat_M11

let ro_M1 = 1/@m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
let ro_M3 = 1/@m.x1.xm3.msky130_fd_pr__nfet_01v8_lvt[gds]
let ro_M5 = 1/@m.x1.xm5.msky130_fd_pr__pfet_01v8_lvt[gds]
let ro_M7 = 1/@m.x1.xm7.msky130_fd_pr__pfet_01v8_lvt[gds]
let ro_M0 = 1/@m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[gds]

print ro_M1
print ro_M3
print ro_M5
print ro_M7
print ro_M0

let gm_M1 = @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm_M3 = @m.x1.xm3.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm_M5 = @m.x1.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm_M7 = @m.x1.xm7.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm_M0 = @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[gm]

print gm_M1
print gm_M3
print gm_M5
print gm_M7
print gm_M0

let gmb_M3 = @m.x1.xm3.msky130_fd_pr__nfet_01v8_lvt[gmbs]
let gmb_M5 = @m.x1.xm5.msky130_fd_pr__pfet_01v8_lvt[gmbs]

print gmb_M3
print gmb_M5


let cgg_M0 = @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[cgg]
print cgg_M0


*CMFB

let x2_vdssat_M0 = @m.x2.xm0.msky130_fd_pr__pfet_01v8_lvt[vdsat]
let x2_vth_M0 = @m.x2.xm0.msky130_fd_pr__pfet_01v8_lvt[vth]

print x2_vdssat_M0
print x2_vth_M0

.endc






.options savecurrents reltol=1e-3 abstol=1e-12 gmin=1e-15
.control
save all

* Operating Point Analysis
op
remzerovec
let cgg_M0 = @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[cgg]
print cgg_M0
write OTA_Telescopic_TB2_STB.raw
set appendwrite

* AC Analysis
ac dec 10 1 5G
remzerovec
write Middlebrook.raw
set appendwrite

* Middlebrook's Method
let tv=-v(vr1)/v(vf1)
let ti=-i(vir1)/i(vif1)
let tmb=(tv*ti - 1)/(tv + ti + 2)

let Av = db(tmb)
meas ac Ao MAX Av
let ABW = Ao-3
meas ac BW WHEN Av=ABW
meas ac UGBW WHEN Av=0

* Phase margin (PM)
let phase_vec= 180/pi*cph(tmb)
meas ac phase FIND phase_vec WHEN frequency=UGBW
let PM = phase+180
print PM

* Gain margin (GM)
meas ac freq180 FIND frequency WHEN phase_vec=-180
meas ac gain FIND Av WHEN frequency=freq180
let GM = 0-gain
print GM

plot Av ylabel 'Magnitude - Middlebrook'
plot phase_vec ylabel 'Phase - Middlebrook'

write Middlebrook_.raw

wrdata STB_Av_ Av
wrdata STB_ph_ phase_vec

*quit

.endc


**** end user architecture code
**.ends

* expanding   symbol:  OTA_Telescopic_core_v2.sym # of pins=8
** sym_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/UNIC-CASS-Aug25/Differential_OTA_Telescopic_IHP/OTA_Telescopic_core_v2.sym
** sch_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/UNIC-CASS-Aug25/Differential_OTA_Telescopic_IHP/OTA_Telescopic_core_v2.sch
.subckt OTA_Telescopic_core_v2 VDD CMFB VOUTP VOUTN VINP VINN VSS IB
*.iopin VDD
*.iopin VSS
*.ipin VINP
*.ipin VINN
*.opin VOUTN
*.opin VOUTP
*.ipin CMFB
*.iopin IB
V2 VB2 VSS 1.5
V3 VB3 VSS 0.7
V4 VB4 VSS 0.49409
V1 VB5 VSS 1.12
* noconn VB2
* noconn VB3
* noconn VB4
* noconn VB5
V5 VB VSS 0.90204
* noconn VB
R1 net1 VOUTP 190 m=1
R2 VOUTN net2 190 m=1
C1 Vo1 net1 0.63p m=1
C2 Vo2 net2 0.63p m=1
XM15 VB55 VB55 VDD VDD sg13_lv_pmos w=1.45u l=0.35u ng=1 m=6
XM17 VB33 VB33 VDD VDD sg13_lv_pmos w=2.05u l=0.35u ng=1 m=1
XM18 VB22 VB33 VDD VDD sg13_lv_pmos w=2.05u l=0.35u ng=1 m=1
XM9 VOUTP Vo1 VDD VDD sg13_lv_pmos w=1.37u l=0.35u ng=1 m=200
XM7 Vx1 VB55 VDD VDD sg13_lv_pmos w=6.85u l=0.7u ng=1 m=30
XM5 Vo1 VB33 Vx1 VDD sg13_lv_pmos w=4.05u l=0.5u ng=1 m=30
XM8 Vx2 VB55 VDD VDD sg13_lv_pmos w=6.85u l=0.7u ng=1 m=30
XM6 Vo2 VB33 Vx2 VDD sg13_lv_pmos w=4.05u l=0.5u ng=1 m=30
XM10 VOUTN Vo2 VDD VDD sg13_lv_pmos w=1.37u l=0.35u ng=1 m=200
XM13 IB IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM14 VB55 IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM16 VB33 IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM19 VB22 VB22 VSS VSS sg13_lv_nmos w=0.5u l=0.8u ng=1 m=1
XM11 VOUTP IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=55
XM0 P CMFB VSS VSS sg13_lv_nmos w=30u l=0.3u ng=9 m=32
XM3 Vo1 VB22 Vy1 VSS sg13_lv_nmos w=1.9u l=0.16u ng=1 m=30
XM1 Vy1 VINP P VSS sg13_lv_nmos w=1.1u l=0.15u ng=1 m=30
XM4 Vo2 VB22 Vy2 VSS sg13_lv_nmos w=1.9u l=0.16u ng=1 m=30
XM2 Vy2 VINN P VSS sg13_lv_nmos w=1.1u l=0.15u ng=1 m=30
XM12 VOUTN IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=55
.ends


* expanding   symbol:  OTA_Telescopic_CMFB2.sym # of pins=7
** sym_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/UNIC-CASS-Aug25/Differential_OTA_Telescopic_IHP/OTA_Telescopic_CMFB2.sym
** sch_path: /foss/designs/Design/xschem/Differential_OTA_Telescopic_IHP/UNIC-CASS-Aug25/Differential_OTA_Telescopic_IHP/OTA_Telescopic_CMFB2.sch
.subckt OTA_Telescopic_CMFB2 VDD VREF VINN VINP IBIAS CMFB VSS
*.iopin VDD
*.iopin VSS
*.opin CMFB
*.ipin VREF
*.iopin IBIAS
*.ipin VINP
*.ipin VINN
XM0 IBIAS IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=8
XM1 V1 IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=24
XM2 V2 IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=24
XM3 CMFB VINP V1 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM4 net1 VREF V1 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM5 net1 VREF V2 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM6 CMFB VINN V2 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM7 net1 net1 VSS VSS sg13_lv_nmos w=30u l=0.3u ng=9 m=6
XM8 CMFB CMFB VSS VSS sg13_lv_nmos w=30u l=0.3u ng=9 m=6
.ends

.GLOBAL GND
.end
