** sch_path: /foss/designs/tb_MUX_4_1.sch
**.subckt tb_MUX_4_1
Vdd4 VDD GND 1.2
Vin2 vinI GND dc 0 ac 0 pulse(0, 1.2, 0, 25p, 25p, 225p, 500p )
Vin1 vinQ GND dc 0 ac 0 pulse(0, 1.2, 125p, 25p, 25p, 225p, 500p )
Vs2 v1 GND 1.2
Vs1 v0 GND 0
Vin3 vinIB GND dc 0 ac 0 pulse(0, 1.2, 250p, 25p, 25p, 225p, 500p )
Vin4 vinQB GND dc 0 ac 0 pulse(0, 1.2, 375p, 25p, 25p, 225p, 500p )
x2 VDD vinI VoutI VoutQ vinQ vinIB VoutIB vinQB VoutQB GND 4to4
x6 v0 VoutI VoutQ VDD Vout v0 v1 VoutIB GND VoutQB MUX_4_1_EN
x1 v0 VoutI VoutQ VDD Vout v1 v1 VoutIB GND VoutQB MUX_4_1_EN
**** begin user architecture code


.param temp=27
.control
save all
tran 0.5p 1.5n

write tran_logic_mux.raw
.endc



.lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends

* expanding   symbol:  4to4.sym # of pins=10
** sym_path: /foss/designs/4to4.sym
** sch_path: /foss/designs/4to4.sch
.subckt 4to4 VDD VINI VOUTI VOUTQ VINQ VINIB VOUTIB VINQB VOUTQB VSS
*.iopin VDD
*.iopin VSS
*.ipin VINI
*.ipin VINQ
*.ipin VINIB
*.ipin VINQB
*.opin VOUTI
*.opin VOUTQ
*.opin VOUTIB
*.opin VOUTQB
x0 VDD net4 VINI VSS inv
x1 VDD net3 VINQ VSS inv
x2 VDD net1 VINIB VSS inv
x3 VDD net2 VINQB VSS inv
x4 VDD VOUTI net4 VSS inv
x5 VDD VOUTQ net3 VSS inv
x6 VDD VOUTIB net1 VSS inv
x7 VDD VOUTQB net2 VSS inv
.ends


* expanding   symbol:  MUX_4_1_EN.sym # of pins=9
** sym_path: /foss/designs/MUX_4_1_EN.sym
** sch_path: /foss/designs/MUX_4_1_EN.sch
.subckt MUX_4_1_EN VEN VINI VINQ VDD VOUT VS[1] VS[0] VINIB VSS VINQB
*.opin VOUT
*.iopin VDD
*.iopin VSS
*.ipin VINI
*.ipin VINQ
*.ipin VINIB
*.ipin VINQB
*.ipin VS[1],VS[0]
*.ipin VEN
x5 VDD net1 net3 VS[1] net2 VSS MUX_2_1
x1 VOUT VEN VENB net3 VDD VSS transmission_gate
x2 VDD VENB VEN VSS inv
x3 VDD VINI net1 VS[0] VINQ VSS MUX_2_1
x4 VDD VINIB net2 VS[0] VINQB VSS MUX_2_1
.ends


* expanding   symbol:  inv.sym # of pins=4
** sym_path: /foss/designs/inv.sym
** sch_path: /foss/designs/inv.sch
.subckt inv VDD VOUT VIN VSS
*.iopin VDD
*.iopin VSS
*.opin VOUT
*.ipin VIN
XM2 VOUT VIN VDD VDD sg13_lv_pmos w=0.15u l=0.13u ng=1 m=2
XM1 VOUT VIN VSS VSS sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
.ends


* expanding   symbol:  MUX_2_1.sym # of pins=6
** sym_path: /foss/designs/MUX_2_1.sym
** sch_path: /foss/designs/MUX_2_1.sch
.subckt MUX_2_1 VDD VINA VOUT VS VINB VSS
*.opin VOUT
*.ipin VINA
*.ipin VINB
*.ipin VS
*.iopin VDD
*.iopin VSS
x1 VOUT net1 VS VINA VDD VSS transmission_gate
x2 VOUT VS net1 VINB VDD VSS transmission_gate
x3 VDD net1 VS VSS inv
.ends


* expanding   symbol:  transmission_gate.sym # of pins=6
** sym_path: /foss/designs/transmission_gate.sym
** sch_path: /foss/designs/transmission_gate.sch
.subckt transmission_gate VOUT VSN VSP VIN VBP VBN
*.iopin VIN
*.iopin VSN
*.iopin VOUT
*.iopin VSP
*.iopin VBN
*.iopin VBP
XM1 VOUT VSN VIN VBN sg13_lv_nmos w=0.15u l=0.13u ng=1 m=1
XM2 VOUT VSP VIN VBP sg13_lv_pmos w=0.15u l=0.13u ng=1 m=2
.ends

.GLOBAL GND
.end
