`default_nettype none   // Prevents implicit net declarations (forces explicit typing)

module uart #(
    parameter NB_DATA      = 32,        // Number of data bits for TX/RX
    parameter NB_STOP      = 16,        // Number of stop bits
    parameter BAUD_RATE    = 19200,     // UART baud rate
    parameter CLK_FREQ     = 45_000_000,// System clock frequency (Hz)
    parameter OVERSAMPLING = 16         // Oversampling factor for sampling RX
)(
    input  wire       clk,        // System clock
    input  wire       i_reset_n,  // Active-low reset
    input  wire       i_rx,       // Serial input line (from external device)
    input  wire [7:0] i_debug2Tx, // Parallel data to transmit (from debug interface)
    input  wire       tx_start,   // Start transmission signal (1 clk pulse)
    output wire       o_tx,       // Serial output line (to external device)
    output wire       o_txDone,   // Transmission completed flag
    output wire       o_rxdone,   // Reception completed flag
    output wire [7:0] o_Rx2debug  // Parallel received data (to debug interface)
);

    // Internal tick signal generated by baudrate_generator
    // Used as a timebase for both RX and TX (oversampled clock)
    wire tick;

    // -------------------------------------------------------------------------
    // Baud rate generator
    // Creates the 'tick' signal based on system clock and configured BAUD_RATE.
    // This tick is used by RX and TX to sample/shift bits at correct intervals.
    // -------------------------------------------------------------------------
    baudrate_generator #(
        .BAUD_RATE    (BAUD_RATE),
        .CLK_FREQ     (CLK_FREQ),
        .OVERSAMPLING (OVERSAMPLING)
    ) baudrate_generator_inst (
        .clk     (clk),        // System clock
        .i_reset (i_reset_n),  // Reset (active-low) passed directly
        .o_tick  (tick)        // Generated tick signal
    );

    // -------------------------------------------------------------------------
    // UART Receiver
    // Samples incoming serial data using 'tick'.
    // Outputs received byte on o_Rx2debug when a frame is complete.
    // -------------------------------------------------------------------------
    uart_rx #(
        .NB_DATA (NB_DATA),
        .NB_STOP (NB_STOP)
    ) uart_rx_inst (
        .clk      (clk),        // System clock
        .i_reset  (i_reset_n),  // Reset (active-low)
        .i_tick   (tick),       // Sampling tick
        .i_data   (i_rx),       // Serial RX line
        .o_data   (o_Rx2debug), // Parallel received data
        .o_rxdone (o_rxdone)    // Reception done pulse
    );

    // -------------------------------------------------------------------------
    // UART Transmitter
    // Shifts out i_debug2Tx serially on o_tx.
    // Controlled by 'tick' to respect baud rate timing.
    // -------------------------------------------------------------------------
    uart_tx #(
        .NB_DATA (NB_DATA),
        .NB_STOP (NB_STOP)
    ) uart_tx_inst (
        .clk        (clk),        // System clock
        .i_reset    (i_reset_n),  // Reset (active-low)
        .i_tick     (tick),       // Transmission tick
        .i_start_tx (tx_start),   // Start transmission
        .i_data     (i_debug2Tx), // Parallel data to send
        .o_txdone   (o_txDone),   // Transmission done pulse
        .o_data     (o_tx)        // Serial TX line
    );

endmodule

`default_nettype wire   // Restore default net type (avoid impacting other files)
