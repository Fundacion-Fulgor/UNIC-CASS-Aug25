** sch_path: /home/designer/shared/UNIC-CASS-Aug25/variable_delay.sch
**.subckt variable_delay VDD_D VIN_D VOUT_D VCONT_D VSS_D
*.iopin VSS_D
*.iopin VDD_D
*.ipin VIN_D
*.opin VOUT_D
*.ipin VCONT_D
XM5 net2 VCONT_D VSS_D VSS_D sg13_lv_nmos w=5u l=0.13u ng=1 m=1
XM6 net1 net3 VDD_D VDD_D sg13_lv_pmos w=5u l=0.13u ng=1 m=1
XM2 VOUT_D VIN_D net1 VDD_D sg13_lv_pmos w=0.88u l=0.13u ng=4 m=1
XM1 VOUT_D VIN_D net2 VSS_D sg13_lv_nmos w=0.4u l=0.13u ng=1 m=1
x1 VDD_D VCONT_D net3 VSS_D inv_1_manual
**.ends

* expanding   symbol:  /home/designer/shared/UNIC-CASS-Aug25/others/inv_1_manual.sym # of pins=4
** sym_path: /home/designer/shared/UNIC-CASS-Aug25/others/inv_1_manual.sym
** sch_path: /home/designer/shared/UNIC-CASS-Aug25/others/inv_1_manual.sch
.subckt inv_1_manual VDD_D A Y VSS_D
*.iopin VDD_D
*.iopin VSS_D
*.iopin A
*.iopin Y
XM1 Y A VSS_D VSS_D sg13_lv_nmos w=10u l=0.13u ng=1 m=1
XM2 Y A VDD_D VDD_D sg13_lv_pmos w=10u l=0.13u ng=1 m=1
.ends

.end
