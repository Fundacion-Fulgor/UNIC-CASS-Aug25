** sch_path: /foss/designs/tb_2x_PI.sch
**.subckt tb_2x_PI
Vin vinQ GND dc 0 ac 0 pulse(0, 1.2, 1n, 1n, 1n, 1n, 4n )
Vin1 vinI GND dc 0 ac 0 pulse(0, 1.2, 0, 1n, 1n, 1n, 4n )
Vdd VDD GND 1.2
XM1 vout vinI GND GND sg13_lv_nmos w=740n l=130n ng=1 m=1
XM2 vout vinI VDD VDD sg13_lv_pmos w=1.48u l=130n ng=1 m=1
XM3 vout vinQ GND GND sg13_lv_nmos w=740n l=130n ng=1 m=1
XM4 vout vinQ VDD VDD sg13_lv_pmos w=1.48u l=130n ng=1 m=1
Vin2 net1 GND dc 0 ac 0 pulse(0, 1.2, 0, 1n, 1n, 1n, 4n )
XM5 voutI net1 GND GND sg13_lv_nmos w=740n l=130n ng=1 m=1
XM6 voutI net1 VDD VDD sg13_lv_pmos w=1.48u l=130n ng=1 m=1
Vin3 net2 GND dc 0 ac 0 pulse(0, 1.2, 1n, 1n, 1n, 1n, 4n )
XM7 voutQ net2 GND GND sg13_lv_nmos w=740n l=130n ng=1 m=1
XM8 voutQ net2 VDD VDD sg13_lv_pmos w=1.48u l=130n ng=1 m=1
**** begin user architecture code


.param temp=27
.control
save all
tran 1p 10n
meas tran tdelay TRIG v(vinI) VAl=0.6 FALl=1 TARG v(vout) VAl=0.6 RISE=1
write tran_logic_not.raw
.endc



.lib cornerMOSlv.lib mos_tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
