** sch_path: /foss/designs/Differential_OTA_Telescopic_IHP/OTA_Telescopic_TB2_OL.sch
**.subckt OTA_Telescopic_TB2_OL
V6 net1 Vcm 0 AC 1
V7 Vcm GND 1.25
V1 VDD GND 1.8
V2 VREF GND dc 0.9 pwl(0 0.8 1u 0.8 1.01u 0.9 0.15m 0.9 0.15m 0)
C1 Vout1 GND 500f m=1
C2 Vout2 GND 500f m=1
R5 net3 Vcm 3k m=1
R6 net4 Vcm 3k m=1
I1 VDD net2 100u
x1 VDD cmfb Vout1 Vout2 net1 Vcm GND net2 OTA_Telescopic_core_v2
x2 VDD VREF Vout1 Vout2 net5 cmfb GND OTA_Telescopic_CMFB2
I2 net5 GND 100u
R1 Vout1 net4 6.72k m=1
R2 Vout2 net3 6.72k m=1
R3 Vcm net4 10G m=1
R4 net1 net3 10G m=1
**** begin user architecture code

** opencircuitdesign pdks install
.lib cornerMOSlv.lib mos_tt
.temp 65



.control
save all
 set color0 = white

* AC simulation
ac dec 1k 1 1T
let Av = db((v(Vout1)-v(Vout2)))
meas ac Ao FIND Av WHEN frequency=10
let ABW = Ao-3
meas ac BW WHEN Av=ABW
meas ac UGBW WHEN Av=0
let phase_vec = 180/pi*cph(v(Vout1)-v(Vout2))

* Phase margin (PM)
meas ac phase FIND phase_vec WHEN frequency=UGBW
let PM = phase+180
print PM

* Gain margin (GM)
meas ac freq180 FIND frequency WHEN phase_vec=-180
meas ac gain FIND Av WHEN frequency=freq180
let GM = 0-gain

*BW in 7 dB
meas ac UGBW7dB WHEN Av=7
meas ac UGBW4dB WHEN Av=4

print GM
plot Av
plot phase_vec

plot db(v(x1.Vo1)-v(x1.Vo2))

write AC_OL.raw

wrdata AvOL_ Av
wrdata PhaseOL_ phase_vec


*DC simulation

op
let vout_dc = v(Vout1)
print vout_dc
write OTA_Telescopic_TB2_OL.raw


reset
noise v(Vout1) V6 dec 100 1 0.5e9 1
setplot noise1
*plot onoise_spectrum
setplot noise2
print onoise_total

.endc




.op

.save all
*OTA
.save @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
.save @m.x1.xm2.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm2.msky130_fd_pr__nfet_01v8_lvt[gm]
.save @m.x1.xm10.msky130_fd_pr__pfet_01v8_lvt[cgg]

.save @m.x1.xm9.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x1.xm9.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x1.xm10.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x1.xm10.msky130_fd_pr__pfet_01v8_lvt[gm]

.save @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[gm]

.save @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[vdssat]


.save @m.x1.xm13.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm13.msky130_fd_pr__nfet_01v8_lvt[gm]
.save @m.x1.xm14.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm15.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x1.xm16.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x1.xm17.msky130_fd_pr__nfet_01v8_lvt[id]

.save @m.x1.xm18.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x1.xm19.msky130_fd_pr__nfet_01v8_lvt[id]

.save @m.x1.xm7.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x1.xm7.msky130_fd_pr__pfet_01v8_lvt[gm]

*CMFB
.save @m.x2.xm0.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm1.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm1.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm2.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm2.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm3.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm3.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm4.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm4.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm5.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
.save @m.x2.xm6.msky130_fd_pr__pfet_01v8_lvt[id]
.save @m.x2.xm6.msky130_fd_pr__pfet_01v8_lvt[gm]

.save @m.x2.xm7.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x2.xm7.msky130_fd_pr__nfet_01v8_lvt[gm]
.save @m.x2.xm8.msky130_fd_pr__nfet_01v8_lvt[id]
.save @m.x2.xm8.msky130_fd_pr__nfet_01v8_lvt[gm]



.control

let vdssat_M1 = @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[vdsat]
let vdssat_M3 = @m.x1.xm3.msky130_fd_pr__nfet_01v8_lvt[vdsat]
let vdssat_M5 = @m.x1.xm5.msky130_fd_pr__pfet_01v8_lvt[vdsat]
let vdssat_M7 = @m.x1.xm7.msky130_fd_pr__pfet_01v8_lvt[vdsat]
let vdssat_M0 = @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[vdsat]

print vdssat_M1
print vdssat_M3
print vdssat_M5
print vdssat_M7
print vdssat_M0

let ro_M1 = 1/@m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[gds]
let ro_M3 = 1/@m.x1.xm3.msky130_fd_pr__nfet_01v8_lvt[gds]
let ro_M5 = 1/@m.x1.xm5.msky130_fd_pr__pfet_01v8_lvt[gds]
let ro_M7 = 1/@m.x1.xm7.msky130_fd_pr__pfet_01v8_lvt[gds]
let ro_M0 = 1/@m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[gds]
let ro_M9 = 1/@m.x1.xm9.msky130_fd_pr__pfet_01v8_lvt[gds]
let ro_M11 = 1/@m.x1.xm11.msky130_fd_pr__nfet_01v8_lvt[gds]

print ro_M1
print ro_M3
print ro_M5
print ro_M7
print ro_M0
print ro_M9
print ro_M11

let gm_M1 = @m.x1.xm1.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm_M3 = @m.x1.xm3.msky130_fd_pr__nfet_01v8_lvt[gm]
let gm_M5 = @m.x1.xm5.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm_M7 = @m.x1.xm7.msky130_fd_pr__pfet_01v8_lvt[gm]
let gm_M0 = @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[gm]

print gm_M1
print gm_M3
print gm_M5
print gm_M7
print gm_M0

let gmb_M3 = @m.x1.xm3.msky130_fd_pr__nfet_01v8_lvt[gmbs]
let gmb_M5 = @m.x1.xm5.msky130_fd_pr__pfet_01v8_lvt[gmbs]

print gmb_M3
print gmb_M5


let cgg_M10 = @m.x1.xm10.msky130_fd_pr__pfet_01v8_lvt[cgg]
print cgg_M10

let cgd_M10 = @m.x1.xm10.msky130_fd_pr__pfet_01v8_lvt[cgd]
print cgd_M10

let cgd_M0 = @m.x1.xm0.msky130_fd_pr__nfet_01v8_lvt[cgd]
print cgd_M0


*CMFB

let x2_vdssat_M0 = @m.x2.xm0.msky130_fd_pr__pfet_01v8_lvt[vdsat]
let x2_vth_M0 = @m.x2.xm0.msky130_fd_pr__pfet_01v8_lvt[vth]

print x2_vdssat_M0
print x2_vth_M0

.endc



**** end user architecture code
**.ends

* expanding   symbol:  OTA_Telescopic_core_v2.sym # of pins=8
** sym_path: /foss/designs/Differential_OTA_Telescopic_IHP/OTA_Telescopic_core_v2.sym
** sch_path: /foss/designs/Differential_OTA_Telescopic_IHP/OTA_Telescopic_core_v2.sch
.subckt OTA_Telescopic_core_v2 VDD CMFB VOUTP VOUTN VINP VINN VSS IB
*.iopin VDD
*.iopin VSS
*.ipin VINP
*.ipin VINN
*.opin VOUTN
*.opin VOUTP
*.ipin CMFB
*.iopin IB
V2 VB2 VSS 1.5
V3 VB3 VSS 0.7
V4 VB4 VSS 0.49409
V1 VB5 VSS 1.12
* noconn VB2
* noconn VB3
* noconn VB4
* noconn VB5
V5 VB VSS 0.90204
* noconn VB
R1 net1 VOUTP 190 m=1
R2 VOUTN net2 190 m=1
C1 Vo1 net1 0.63p m=1
C2 Vo2 net2 0.63p m=1
XM15 VB55 VB55 VDD VDD sg13_lv_pmos w=1.45u l=0.35u ng=1 m=6
XM17 VB33 VB33 VDD VDD sg13_lv_pmos w=2.05u l=0.35u ng=1 m=1
XM18 VB22 VB33 VDD VDD sg13_lv_pmos w=2.05u l=0.35u ng=1 m=1
XM9 VOUTP Vo1 VDD VDD sg13_lv_pmos w=1.37u l=0.35u ng=1 m=200
XM7 Vx1 VB55 VDD VDD sg13_lv_pmos w=6.85u l=0.7u ng=1 m=30
XM5 Vo1 VB33 Vx1 VDD sg13_lv_pmos w=4.05u l=0.5u ng=1 m=30
XM8 Vx2 VB55 VDD VDD sg13_lv_pmos w=6.85u l=0.7u ng=1 m=30
XM6 Vo2 VB33 Vx2 VDD sg13_lv_pmos w=4.05u l=0.5u ng=1 m=30
XM10 VOUTN Vo2 VDD VDD sg13_lv_pmos w=1.37u l=0.35u ng=1 m=200
XM13 IB IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM14 VB55 IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM16 VB33 IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=1
XM19 VB22 VB22 VSS VSS sg13_lv_nmos w=0.5u l=0.8u ng=1 m=1
XM11 VOUTP IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=55
XM0 P CMFB VSS VSS sg13_lv_nmos w=57u l=0.3u ng=12 m=16
XM3 Vo1 VB22 Vy1 VSS sg13_lv_nmos w=1.9u l=0.16u ng=1 m=30
XM1 Vy1 VINP P VSS sg13_lv_nmos w=1.1u l=0.15u ng=1 m=30
XM4 Vo2 VB22 Vy2 VSS sg13_lv_nmos w=1.9u l=0.16u ng=1 m=30
XM2 Vy2 VINN P VSS sg13_lv_nmos w=1.1u l=0.15u ng=1 m=30
XM12 VOUTN IB VSS VSS sg13_lv_nmos w=4.8u l=1.06u ng=1 m=55
.ends


* expanding   symbol:  OTA_Telescopic_CMFB2.sym # of pins=7
** sym_path: /foss/designs/Differential_OTA_Telescopic_IHP/OTA_Telescopic_CMFB2.sym
** sch_path: /foss/designs/Differential_OTA_Telescopic_IHP/OTA_Telescopic_CMFB2.sch
.subckt OTA_Telescopic_CMFB2 VDD VREF VINN VINP IBIAS CMFB VSS
*.iopin VDD
*.iopin VSS
*.opin CMFB
*.ipin VREF
*.iopin IBIAS
*.ipin VINP
*.ipin VINN
XM0 IBIAS IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=8
XM1 V1 IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=24
XM2 V2 IBIAS VDD VDD sg13_lv_pmos w=6u l=0.7u ng=6 m=24
XM3 CMFB VINP V1 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM4 net1 VREF V1 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM5 net1 VREF V2 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM6 CMFB VINN V2 VDD sg13_lv_pmos w=9u l=0.35u ng=7 m=4
XM7 net1 net1 VSS VSS sg13_lv_nmos w=57u l=0.3u ng=50 m=4
XM8 CMFB CMFB VSS VSS sg13_lv_nmos w=57u l=0.3u ng=50 m=4
.ends

.GLOBAL GND
.end
